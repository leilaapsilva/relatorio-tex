library verilog;
use verilog.vl_types.all;
entity verilogmerda_vlg_vec_tst is
end verilogmerda_vlg_vec_tst;
