library verilog;
use verilog.vl_types.all;
entity Cenario2_vlg_check_tst is
    port(
        LEDR            : in     vl_logic_vector(1 downto 1);
        sampler_rx      : in     vl_logic
    );
end Cenario2_vlg_check_tst;
