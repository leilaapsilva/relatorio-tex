library verilog;
use verilog.vl_types.all;
entity LLDX_vlg_vec_tst is
end LLDX_vlg_vec_tst;
