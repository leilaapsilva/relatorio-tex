library verilog;
use verilog.vl_types.all;
entity Cenario2_vlg_vec_tst is
end Cenario2_vlg_vec_tst;
