library verilog;
use verilog.vl_types.all;
entity asd123_vlg_vec_tst is
end asd123_vlg_vec_tst;
